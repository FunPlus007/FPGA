// exp 10 mod 24 counter
// 奇怪的要求不知道了 后面在看这个沙雕

module counter_mod24();

endmodule